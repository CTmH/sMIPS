`timescale 1ns / 1ps
module bus(
           input wire sck,
           input wire rst
)
